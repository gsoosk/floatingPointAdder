module Adder(input[24:0] N1, N2, output[24:0] Answer);
  assign Answer = N1 + N2;
endmodule
