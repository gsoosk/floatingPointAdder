module TB();
  //4.56
  reg [31:0] Ain = 32'b01000000100100011110101110000101;
  //-2.12
  reg [31:0] Bin = 32'b11000000000001111010111000010100;
  //ans : 2.14
  
  
  //reg [31:0] Ain = 32'b01000011000010000101011100001010;
  //reg [31:0] Bin = 32'b11000010010110101010111000010100;
  
  //2.5
  //reg [31:0] Ain = 32'b01000000001000000000000000000000 ;
  //1.25
  //reg [31:0] Bin = 32'b00111111101000000000000000000000;
  //ans : 3.75 : 01000000011100000000000000000000
  
  //-2.55
  //reg [31:0] Ain = 32'b11000000001000110011001100110011 ;
  //-4.76
  //reg [31:0] Bin = 32'b11000000100110000101000111101100;
  //ans : -7.31 : 11000000111010011110101110000101




  
  
  
  reg start = 0;
  reg clk=0;
  reg rst = 1 ;
  wire done;
  wire [31:0] Ans;
  
  
  
  floatingPointAdder uut( Ain, Bin, clk, rst, start , done, Ans);
  initial repeat(270) #12 clk=~clk;
  initial begin
    #30 rst=0;
    #50 start=1;
    #70 start=0;
    
  end  
endmodule
