module Adder(input[25:0] N1, N2, output[25:0] Answer);
  assign Answer = N1 + N2;
endmodule
